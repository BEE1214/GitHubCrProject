--=================================--
--=-Project: ProjectName-------------=--
--=-Author: Adam Dvorsky----------=--
--=-Date: date -------------=--
--=================================--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- use IEEE.NUMERIC_STD.ALL;

entity $argv[1] is
  port (
    CLK : in std_logic;
  ) ;
end $argv[1];

